`define NBIT 8
`define KERNEL_SIZE 3
`define NBIT_SOBEL 16
//tb params
`define NUM_TESTS 5
`define FRAC_BITS 10