`define NBIT 8
`define KERNEL_SIZE 3

//tb params
`define NUM_TESTS 100
`define FRAC_BITS 10