`define NBIT 8
`define KERNEL_SIZE 3
`define NBIT_SOBEL 16

//ARCTANG LUT SIZE
`define LUT_ATAN_SIZE 1024
//tb params
`define NUM_TESTS 5
`define FRAC_BITS 10